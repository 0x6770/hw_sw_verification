package pkg;
  `include "transaction.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "test.sv"
  `include "environment.sv"
endpackage
