import pkg::*;

module environment;
  AHB_monitor monitor;
  AHB_driver driver;
  AHB_scoreboard scoreboard;
endmodule
