module test #(
    parameter byte GPIO_DATA_ADDR = 8'h00,
    parameter byte GPIO_DIR_ADDR  = 8'h04
) ();
endmodule
