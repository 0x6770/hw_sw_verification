package pkg;
  `include "transaction.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "generator.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
endpackage
