package pkg;
  // `include "transaction.sv"
  // `include "driver.sv"
  // `include "monitor.sv"
  // `include "generator.sv"
  // `include "scoreboard.sv"
  `include "environment.sv"
  // `include "ahb_pkg.sv"
  // `include "ahb_gpio.sv"
endpackage
